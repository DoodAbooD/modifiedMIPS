module test(in, out);
    

endmodule